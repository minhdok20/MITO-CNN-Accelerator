//`timescale 1ns / 1ps

//module CONTROLLER #(parameter ) 
//                   ();
                   
    
    
//endmodule
